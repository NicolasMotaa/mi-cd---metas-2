module and8bits (S, A, B);

	output [7:0] S;
	input  [7:0] A;
	input  [7:0] B;

	and And0 (S[0], A[0], B[0]);
	and And1 (S[1], A[1], B[1]);
	and And2 (S[2], A[2], B[2]);
	and And3 (S[3], A[3], B[3]);
	and And4 (S[4], A[4], B[4]);
	and And5 (S[5], A[5], B[5]);
	and And6 (S[6], A[6], B[6]);
	and And7 (S[7], A[7], B[7]);

endmodule
